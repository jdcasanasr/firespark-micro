// Fetch stage parameters.
`define ICACHE_DEPTH 128