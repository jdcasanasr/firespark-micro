`define XLEN 32